import common::*;
module video(
    input rst_n,
    input clk28,

    input machine_t machine,
    input [2:0] border,
    input up_en,

    output reg [2:0] r,
    output reg [2:0] g,
    output reg [1:0] b,
    output reg vsync,
    output reg hsync,
    output reg csync,

    output read_req,
    output read_req_is_up,
    output [14:0] read_req_addr,
    input read_req_ack,
    input read_data_valid,
    input [7:0] read_data,

    output contention,
    output reg even_line,
    output port_ff_active,
    output [7:0] port_ff_data,

    output [8:0] hc_out,
    output [8:0] vc_out,
    output clk14,
    output clk7,
    output clk35,
    output ck14,
    output ck7,
    output ck35,
    output clk25hz,
    output clk12_5hz,
    output clk6_25hz,
    output clk3_125hz,
    output clk1_5625hz,
    input [5:0] timex_mode,
    output ext_palette
);

reg  [8:0] vc;
reg  [10:0] hc0;
wire [8:0] hc = hc0[10:2];
assign vc_out = vc;
assign hc_out = hc;

assign clk14 = hc0[0];
assign clk7 = hc0[1];
assign clk35 = hc0[2];
assign ck14 = hc0[0];
assign ck7 = hc0[0] & hc0[1];
assign ck35 = hc0[0] & hc0[1] & hc0[2];

reg [4:0] blink_cnt;
assign clk25hz = blink_cnt[0];
assign clk12_5hz = blink_cnt[1];
assign clk6_25hz = blink_cnt[2];
assign clk3_125hz = blink_cnt[3];
assign clk1_5625hz = blink_cnt[4];


/* SYNC SIGNALS */
localparam H_AREA         = 256;
localparam V_AREA         = 192;
localparam SCREEN_DELAY   = 13;

localparam H_LBORDER_S48  = 54 - SCREEN_DELAY;
localparam H_RBORDER_S48  = 53 + SCREEN_DELAY;
localparam H_BLANK1_S48   = 12;
localparam H_SYNC_S48     = 33;
localparam H_BLANK2_S48   = 40;
localparam H_TOTAL_S48    = H_AREA + H_RBORDER_S48 + H_BLANK1_S48 + H_SYNC_S48 + H_BLANK2_S48 + H_LBORDER_S48;
localparam V_BBORDER_S48  = 56;
localparam V_SYNC_S48     = 8;
localparam V_TBORDER_S48  = 56;
localparam V_TOTAL_S48    = V_AREA + V_BBORDER_S48 + V_SYNC_S48 + V_TBORDER_S48;

localparam H_LBORDER_S128 = 54 - SCREEN_DELAY;
localparam H_RBORDER_S128 = 53 + SCREEN_DELAY;
localparam H_BLANK1_S128  = 16;
localparam H_SYNC_S128    = 33;
localparam H_BLANK2_S128  = 44;
localparam H_TOTAL_S128   = H_AREA + H_RBORDER_S128 + H_BLANK1_S128 + H_SYNC_S128 + H_BLANK2_S128 + H_LBORDER_S128;
localparam V_BBORDER_S128 = 55;
localparam V_SYNC_S128    = 8;
localparam V_TBORDER_S128 = 56;
localparam V_TOTAL_S128   = V_AREA + V_BBORDER_S128 + V_SYNC_S128 + V_TBORDER_S128;

localparam H_LBORDER_PENT = 54 - SCREEN_DELAY;
localparam H_RBORDER_PENT = 53 + SCREEN_DELAY;
localparam H_BLANK1_PENT  = 12;
localparam H_SYNC_PENT    = 33;
localparam H_BLANK2_PENT  = 40;
localparam H_TOTAL_PENT   = H_AREA + H_RBORDER_PENT + H_BLANK1_PENT + H_SYNC_PENT + H_BLANK2_PENT + H_LBORDER_PENT;
localparam V_BBORDER_PENT = 56;
localparam V_SYNC_PENT    = 8;
localparam V_TBORDER_PENT = 64;
localparam V_TOTAL_PENT   = V_AREA + V_BBORDER_PENT + V_SYNC_PENT + V_TBORDER_PENT;

wire hc0_reset =
    (machine == MACHINE_S48)?
        hc0 == (H_TOTAL_S48<<2) - 1'b1 :
    (machine == MACHINE_S128 || machine == MACHINE_S3)?
        hc0 == (H_TOTAL_S128<<2) - 1'b1 :
    // Pentagon
        hc0 == (H_TOTAL_PENT<<2) - 1'b1 ;
wire vc_reset =
    (machine == MACHINE_S48)?
        vc == V_TOTAL_S48 - 1'b1:
    (machine == MACHINE_S128 || machine == MACHINE_S3)?
        vc == V_TOTAL_S128 - 1'b1 :
    // Pentagon
        vc == V_TOTAL_PENT - 1'b1 ;
wire hsync0 =
    (machine == MACHINE_S48)?
        (hc >= (H_AREA + H_RBORDER_S48 + H_BLANK1_S48)) && (hc < (H_AREA + H_RBORDER_S48 + H_BLANK1_S48 + H_SYNC_S48)) :
    (machine == MACHINE_S128 || machine == MACHINE_S3)?
        (hc >= (H_AREA + H_RBORDER_S128 + H_BLANK1_S128)) && (hc < (H_AREA + H_RBORDER_S128 + H_BLANK1_S128 + H_SYNC_S128)) :
    // Pentagon
        (hc >= (H_AREA + H_RBORDER_PENT + H_BLANK1_PENT)) && (hc < (H_AREA + H_RBORDER_PENT + H_BLANK1_PENT + H_SYNC_PENT)) ;
wire vsync0 =
    (machine == MACHINE_S48)?
        (vc >= (V_AREA + V_BBORDER_S48)) && (vc < (V_AREA + V_BBORDER_S48 + V_SYNC_S48)) :
    (machine == MACHINE_S128 || machine == MACHINE_S3)?
        (vc >= (V_AREA + V_BBORDER_S128)) && (vc < (V_AREA + V_BBORDER_S128 + V_SYNC_S128)) :
    // Pentagon
        (vc >= (V_AREA + V_BBORDER_PENT)) && (vc < (V_AREA + V_BBORDER_PENT + V_SYNC_PENT)) ;
wire blank =
    (machine == MACHINE_S48)?
        ((vc >= (V_AREA + V_BBORDER_S48)) && (vc < (V_AREA + V_BBORDER_S48 + V_SYNC_S48))) ||
            ((hc >= (H_AREA + H_RBORDER_S48)) &&
             (hc <  (H_AREA + H_RBORDER_S48 + H_BLANK1_S48 + H_SYNC_S48 + H_BLANK2_S48))) :
    (machine == MACHINE_S128 || machine == MACHINE_S3)?
        ((vc >= (V_AREA + V_BBORDER_S128)) && (vc < (V_AREA + V_BBORDER_S128 + V_SYNC_S128))) ||
            ((hc >= (H_AREA + H_RBORDER_S128)) &&
             (hc <  (H_AREA + H_RBORDER_S128 + H_BLANK1_S128 + H_SYNC_S128 + H_BLANK2_S128))) :
    // Pentagon
        ((vc >= (V_AREA + V_BBORDER_PENT)) && (vc < (V_AREA + V_BBORDER_PENT + V_SYNC_PENT))) ||
            ((hc >= (H_AREA + H_RBORDER_PENT)) &&
             (hc <  (H_AREA + H_RBORDER_PENT + H_BLANK1_PENT + H_SYNC_PENT + H_BLANK2_PENT))) ;

always @(posedge clk28 or negedge rst_n) begin
    if (!rst_n) begin
        hc0 <= 0;
        vc <= 0;
    end
    else if (hc0_reset) begin
        hc0 <= 0;
        if (vc_reset) begin
            vc <= 0;
        end
        else begin
            vc <= vc + 1'b1;
        end
    end
    else begin
        hc0 <= hc0 + 1'b1;
    end
end

wire blink = blink_cnt[$bits(blink_cnt)-1];
always @(posedge clk28 or negedge rst_n) begin
    if (!rst_n)
        blink_cnt <= 0;
    else if (hc0_reset && vc_reset)
        blink_cnt <= blink_cnt + 1'b1;
end

reg hsync0_delayed;
always @(posedge clk28)
    hsync0_delayed <= hsync0;
always @(posedge clk28 or negedge rst_n) begin
    if (!rst_n)
        even_line <= 0;
    else if (hsync0 && !hsync0_delayed)
        even_line <= ~even_line;
end


/* SCREEN CONTROLLER */

wire timex_page = timex_mode[0] & ~timex_mode[2] & ~timex_mode[1];
wire timex_hi_col = timex_mode[1];
wire timex_hi_res = timex_mode[2] & ~timex_mode[0]; // must be set together with [1]

// 4colors modes need all HiResColors bits, so the forbidden combinations are used
wire CGA_mode4col = timex_mode[2] & timex_mode[1] & timex_mode[0];
wire BiPlanes_mode4col = ~timex_mode[2] & timex_mode[1] & timex_mode[0]; // Dual Playfield mode
wire CGA_mode16col = up_en & timex_mode[3] & ~timex_mode[2] & ~timex_mode[1];// & ~timex_mode[0];

wire screen_show = (vc < V_AREA) && (hc0 >= (SCREEN_DELAY<<2) - 1) && (hc0 < ((H_AREA + SCREEN_DELAY)<<2) - 1);
wire screen_update = hc0[4:0] == 5'b10011;
wire border_update = (hc0[4:0] == 5'b10011) || (machine == MACHINE_PENT && ck7);
wire bitmap_shift = hc0[1:0] == 2'b11 && ! (CGA_mode16col || BiPlanes_mode4col)  // 128 cols
  || hc0[2:0] == 3'b011               // 256 cols
  || timex_hi_res && hc0[0] == 1'b1;  // 512 cols
wire next_addr = hc0[4:0] == 5'b10001;

reg screen_read;
always @(posedge clk28)
    screen_read <= (vc < V_AREA) && (hc0 > 17) && (hc0 < (H_AREA<<2) + 17);

reg [7:0] vaddr;
reg [7:3] haddr;
always @(posedge clk28 or negedge rst_n) begin
    if (!rst_n) begin
        vaddr <= 0;
        haddr <= 0;
    end
    else if (next_addr) begin
        vaddr <= vc[7:0];
        haddr <= hc[7:3];
    end
end

reg [7:0] bitmap, attr, bitmap_next, attr_next, bitmap_odd, bitmap_odd_next;
reg [7:0] up_ink, up_paper, up_ink_next, up_paper_next;
reg [7:0] up_col11, up_col01; // second ink, second paper in 4 in 16 color modes
reg colors01and11;

reg [1:0] read_step, read_step_cur;
assign read_req = 1'b1; // just to simplify logic
// TIMEX MULTICOLOR atribute address / HiRes OddColumn, CGA 4 and 16 color modes:
wire read_2nd_page = timex_hi_col | CGA_mode16col; //| CGA_mode4col | BiPlanes_mode4col);
assign read_req_addr =
    (read_step == 2'd3)? { attr_next[7:6], 1'b1, attr_next[5:3] } :
    ((read_step == 2'd2)
              && up_en)? { attr_next[7:6], 1'b0, attr_next[2:0] } :
    (read_step == 2'd1)? { 1'b1, timex_page, vaddr[7:6], vaddr[2:0], vaddr[5:3], haddr[7:3] } :
    (read_2nd_page && read_step == 2'd0)?
                         { 2'b11, vaddr[7:6], vaddr[2:0], vaddr[5:3], haddr[7:3] } :
                         { 1'b1, timex_page, 3'b110, vaddr[7:3], haddr[7:3] } ;

assign read_req_is_up = (read_step == 2'd2 && up_en) || (read_step == 2'd3);
assign ext_palette = up_en | CGA_mode4col | CGA_mode16col | BiPlanes_mode4col;

always @(posedge clk28 or negedge rst_n) begin
    if (!rst_n) begin
        read_step <= 0;
        read_step_cur <= 0;
        attr_next <= 0;
        bitmap_next <= 0;
        up_ink_next <= 0;
        up_paper_next <= 0;
        bitmap_odd_next <= 0;
        colors01and11 <= 0;
    end
    else begin
        if (next_addr)
            read_step <= 0;
        else if (read_req_ack && !(up_en | CGA_mode4col | BiPlanes_mode4col) && read_step[0])
            read_step <= 0;
        else if (read_req_ack && !(up_en) && read_step[1])
            read_step <= 0;
        else if (read_req_ack)
            read_step <= read_step + 1'd1;

        if (read_req_ack)
            read_step_cur <= read_step;

        if (read_data_valid && read_step_cur == 2'd0 && screen_read) begin
            if (~read_2nd_page | ~(timex_hi_res | CGA_mode4col | CGA_mode16col | BiPlanes_mode4col))
                attr_next <= read_data;  // in step "0" regular ZX or Timex HiCol attributes are read
            else if (read_2nd_page) begin
                bitmap_odd_next <= read_data;
                if (timex_hi_res)
                    attr_next <= {1'b0, up_en, ~timex_mode[5:3], timex_mode[5:3]};
                else if (up_en & (CGA_mode4col | CGA_mode16col | BiPlanes_mode4col)) begin
                    colors01and11 <= haddr[3] & ~CGA_mode4col;
                    // just to allow proper ULA+ reading "zones" for colors
                    attr_next <= { ~vaddr[7:6], vaddr[5:4], 
                            CGA_mode4col ? vaddr[3] : haddr[3],
                            vaddr[5:4],
                            CGA_mode4col ? vaddr[3] : haddr[3]};
                end
            end
        end
        else if (!screen_read && hc0[0]) begin
            // timex HiRes keeps paper color on border.
            if (~timex_hi_res)
                attr_next <= {1'b0, up_en, ~timex_mode[5:3], ~timex_mode[5:3]};
            if (~up_en)
                up_paper_next <= color16_256({1'b0, border[2:0]});
            bitmap_odd_next <= 0;
        end

        if (read_data_valid && read_step_cur == 2'd1 && screen_read)
            bitmap_next <= read_data;
        else if (!screen_read && hc0[0]) begin
            bitmap_next <= 0;
        end

        if (read_data_valid && read_step_cur == 2'd2) begin
            // step 2 is either ULA+ ink read from pallette
            // either CGA4 or DualPlayField attributes read
            if (!up_en && screen_read) begin 
                up_ink_next <= color16_256(read_data[3:0]);
                up_paper_next <= color16_256(read_data[7:4]);
                colors01and11 <= 1'b0;
            end
            else
                up_ink_next <= read_data;
        end
        if (read_data_valid && read_step_cur == 2'd3)
            up_paper_next <= read_data;
    end
end

always @(posedge clk28 or negedge rst_n) begin
    if (!rst_n) begin
        attr <= 0;
        bitmap <= 0;
        bitmap_odd <= 0;
        up_ink <= 0;
        up_paper <= 0;
        up_col11 <= 0;
        up_col01 <= 0;
    end
    else begin
        if (screen_show && screen_update) begin
            attr <= attr_next;
        end
        else if (!screen_show && border_update) begin
            attr <= {2'b00, border[2:0], border[2:0]};
            // in CGA-style modes, the up_paper_next arleady contains proper border color
            // it also works in all ULA+ cases
            if (ext_palette)
                up_paper = up_paper_next;
        end

        if (screen_update) begin
            bitmap <= bitmap_next;
            bitmap_odd <= bitmap_odd_next;
        end
        else if (bitmap_shift)
            if (CGA_mode4col | BiPlanes_mode4col) begin
                bitmap <= {bitmap[5:0], bitmap_odd[7:6]};
                bitmap_odd <= {bitmap_odd[5:0], 2'b00};
            end
            else if (CGA_mode16col) begin
                bitmap <= {bitmap[3:0], bitmap_odd[7:4]};
                bitmap_odd <= {bitmap_odd[3:0], 4'b0000};
            end
            else begin
                bitmap <= {bitmap[6:0], bitmap_odd[7]};
                bitmap_odd <= {bitmap_odd[6:0], 1'b0};
            end
        if (screen_update)
            if (colors01and11) begin
                up_col11 <= up_ink_next;
                up_col01 <= up_paper_next;
            end
            else begin
                up_ink <= up_ink_next;
                up_paper <= up_paper_next;
            end
    end
end

/* ATTRIBUTE PORT */
wire port_ff_attr = (machine == MACHINE_PENT) || hc[3:1] == 3'h6 || hc[3:1] == 3'h0;
wire port_ff_bitmap = (hc[3] && hc[1]);
assign port_ff_active = screen_read && (port_ff_attr || port_ff_bitmap);
assign port_ff_data =
    port_ff_attr? attr_next :
    port_ff_bitmap? bitmap_next :
    8'hFF;

assign contention = (vc < V_AREA) && (hc < H_AREA) && (hc[2] || hc[3]);

function [7:0] color16_256; input [4:0] in;
    color16_256 = {in[2], in[2] | in[3], 1'b0, // G
                   in[1] | in[3], in[1], 1'b0, // R
                   in[0], in[0]};      // B
endfunction

/* RGBS OUTPUT */
wire second_playfield = BiPlanes_mode4col && bitmap[7:6] == 2'b11;
wire pixel = second_playfield ?
        bitmap_odd[7] :
        bitmap[7];
wire second_colpair_selector = 
    (CGA_mode16col | BiPlanes_mode4col | CGA_mode4col) ?
        ( second_playfield ?
            bitmap_odd[6] :
            bitmap[6]
        ) :
        1'b0;
// in 16Col mode, 12 colors is direct, rest is from ULAPlus
wire CGA_mode16col_direct = screen_show && CGA_mode16col & (~(bitmap[7] ^ bitmap[4]) | bitmap[5]);

always @* begin
    if (blank)
        {g, r, b} = 0;
    else if (CGA_mode16col_direct) begin
        {g, r, b} = color16_256(bitmap[7:4]);
    end
    else if (ext_palette & ~second_colpair_selector & ~second_playfield) begin
        g = pixel? up_ink[7:5] : up_paper[7:5];
        r = pixel? up_ink[4:2] : up_paper[4:2];
        b = pixel? up_ink[1:0] : up_paper[1:0];
    end
    else if (second_colpair_selector & CGA_mode16col | second_playfield & ~second_colpair_selector) begin
        g = pixel? up_col11[7:5] : up_col01[7:5];
        r = pixel? up_col11[4:2] : up_col01[4:2];
        b = pixel? up_col11[1:0] : up_col01[1:0];
    end
    else if (second_colpair_selector && (BiPlanes_mode4col | CGA_mode4col))
            // for 11 choose additional Timex color, for 01 choose second page point colors + border + combined
            {g, r, b} = 
                (~pixel) ? color16_256({second_playfield, border[2:0]}) :
                        color16_256 ({~second_playfield, timex_mode[5:3]});
    else begin
        {g[2], r[2], b[1]} = (pixel ^ (attr[7] & blink))? attr[2:0] : attr[5:3];
        {g[1], r[1], b[0]} = ((g[2] | r[2] | b[1]) & attr[6])? 3'b111 : 3'b000;
        {g[0], r[0]} = 2'b00;
    end
end

always @(posedge clk28) begin
    csync = ~(vsync0 ^ hsync0);
    vsync = vsync0;
    hsync = hsync0;
end


endmodule
